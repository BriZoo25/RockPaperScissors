module ScoreSeven (input [3:0]i, output reg [6:0]o);
	
	always@(*)
		begin
			case(i)
				4'b0000: o = 7'b0000001;//0
				4'b0001: o = 7'b1001111;//1
				4'b0010: o = 7'b0010010;//2
				4'b0011: o = 7'b0000110;//3
				4'b0100: o = 7'b1001100;//4
				4'b0101: o = 7'b0100100;//5
				4'b0110: o = 7'b0100000;//6
				4'b0111: o = 7'b0001111;//7
				4'b1000: o = 7'b0000000;//8
				4'b1001: o = 7'b0001100;//9
				
				
				default: o = 7'b1111111;
			endcase
		end
endmodule 